library verilog;
use verilog.vl_types.all;
entity cnt3reset4_vlg_vec_tst is
end cnt3reset4_vlg_vec_tst;
