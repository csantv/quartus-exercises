library verilog;
use verilog.vl_types.all;
entity cnt5reset23_vlg_vec_tst is
end cnt5reset23_vlg_vec_tst;
