library verilog;
use verilog.vl_types.all;
entity lab2p2_vlg_check_tst is
    port(
        COMESTIBLES     : in     vl_logic;
        MEDICINAS       : in     vl_logic;
        TECNOLOGIA      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab2p2_vlg_check_tst;
