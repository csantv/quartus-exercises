library verilog;
use verilog.vl_types.all;
entity lab2p2_vlg_vec_tst is
end lab2p2_vlg_vec_tst;
