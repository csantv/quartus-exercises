library verilog;
use verilog.vl_types.all;
entity cnt3reset4_vlg_check_tst is
    port(
        Out0            : in     vl_logic;
        Out1            : in     vl_logic;
        Out2            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end cnt3reset4_vlg_check_tst;
